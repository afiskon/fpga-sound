/* vim: set ai et ts=4 sw=4: */
`default_nettype none

module sine_sig(input logic clk, output logic [0:7] sig);
    logic [0:7] counter;

    sawtooth_sig st_sig(clk, counter);

    always_ff @(posedge clk)
    begin
        case (counter)

            8'b00000000: sig <= 8'b01111111;
            8'b00000001: sig <= 8'b10000010;
            8'b00000010: sig <= 8'b10000101;
            8'b00000011: sig <= 8'b10001000;
            8'b00000100: sig <= 8'b10001011;
            8'b00000101: sig <= 8'b10001110;
            8'b00000110: sig <= 8'b10010001;
            8'b00000111: sig <= 8'b10010100;
            8'b00001000: sig <= 8'b10010111;
            8'b00001001: sig <= 8'b10011010;
            8'b00001010: sig <= 8'b10011101;
            8'b00001011: sig <= 8'b10100000;
            8'b00001100: sig <= 8'b10100011;
            8'b00001101: sig <= 8'b10100110;
            8'b00001110: sig <= 8'b10101001;
            8'b00001111: sig <= 8'b10101100;
            8'b00010000: sig <= 8'b10101111;
            8'b00010001: sig <= 8'b10110010;
            8'b00010010: sig <= 8'b10110101;
            8'b00010011: sig <= 8'b10111000;
            8'b00010100: sig <= 8'b10111010;
            8'b00010101: sig <= 8'b10111101;
            8'b00010110: sig <= 8'b11000000;
            8'b00010111: sig <= 8'b11000010;
            8'b00011000: sig <= 8'b11000101;
            8'b00011001: sig <= 8'b11001000;
            8'b00011010: sig <= 8'b11001010;
            8'b00011011: sig <= 8'b11001101;
            8'b00011100: sig <= 8'b11001111;
            8'b00011101: sig <= 8'b11010001;
            8'b00011110: sig <= 8'b11010100;
            8'b00011111: sig <= 8'b11010110;
            8'b00100000: sig <= 8'b11011000;
            8'b00100001: sig <= 8'b11011010;
            8'b00100010: sig <= 8'b11011101;
            8'b00100011: sig <= 8'b11011111;
            8'b00100100: sig <= 8'b11100001;
            8'b00100101: sig <= 8'b11100011;
            8'b00100110: sig <= 8'b11100101;
            8'b00100111: sig <= 8'b11100110;
            8'b00101000: sig <= 8'b11101000;
            8'b00101001: sig <= 8'b11101010;
            8'b00101010: sig <= 8'b11101011;
            8'b00101011: sig <= 8'b11101101;
            8'b00101100: sig <= 8'b11101111;
            8'b00101101: sig <= 8'b11110000;
            8'b00101110: sig <= 8'b11110001;
            8'b00101111: sig <= 8'b11110011;
            8'b00110000: sig <= 8'b11110100;
            8'b00110001: sig <= 8'b11110101;
            8'b00110010: sig <= 8'b11110110;
            8'b00110011: sig <= 8'b11110111;
            8'b00110100: sig <= 8'b11111000;
            8'b00110101: sig <= 8'b11111001;
            8'b00110110: sig <= 8'b11111010;
            8'b00110111: sig <= 8'b11111010;
            8'b00111000: sig <= 8'b11111011;
            8'b00111001: sig <= 8'b11111100;
            8'b00111010: sig <= 8'b11111100;
            8'b00111011: sig <= 8'b11111101;
            8'b00111100: sig <= 8'b11111101;
            8'b00111101: sig <= 8'b11111101;
            8'b00111110: sig <= 8'b11111101;
            8'b00111111: sig <= 8'b11111101;
            8'b01000000: sig <= 8'b11111110;
            8'b01000001: sig <= 8'b11111101;
            8'b01000010: sig <= 8'b11111101;
            8'b01000011: sig <= 8'b11111101;
            8'b01000100: sig <= 8'b11111101;
            8'b01000101: sig <= 8'b11111101;
            8'b01000110: sig <= 8'b11111100;
            8'b01000111: sig <= 8'b11111100;
            8'b01001000: sig <= 8'b11111011;
            8'b01001001: sig <= 8'b11111010;
            8'b01001010: sig <= 8'b11111010;
            8'b01001011: sig <= 8'b11111001;
            8'b01001100: sig <= 8'b11111000;
            8'b01001101: sig <= 8'b11110111;
            8'b01001110: sig <= 8'b11110110;
            8'b01001111: sig <= 8'b11110101;
            8'b01010000: sig <= 8'b11110100;
            8'b01010001: sig <= 8'b11110011;
            8'b01010010: sig <= 8'b11110001;
            8'b01010011: sig <= 8'b11110000;
            8'b01010100: sig <= 8'b11101111;
            8'b01010101: sig <= 8'b11101101;
            8'b01010110: sig <= 8'b11101011;
            8'b01010111: sig <= 8'b11101010;
            8'b01011000: sig <= 8'b11101000;
            8'b01011001: sig <= 8'b11100110;
            8'b01011010: sig <= 8'b11100101;
            8'b01011011: sig <= 8'b11100011;
            8'b01011100: sig <= 8'b11100001;
            8'b01011101: sig <= 8'b11011111;
            8'b01011110: sig <= 8'b11011101;
            8'b01011111: sig <= 8'b11011010;
            8'b01100000: sig <= 8'b11011000;
            8'b01100001: sig <= 8'b11010110;
            8'b01100010: sig <= 8'b11010100;
            8'b01100011: sig <= 8'b11010001;
            8'b01100100: sig <= 8'b11001111;
            8'b01100101: sig <= 8'b11001101;
            8'b01100110: sig <= 8'b11001010;
            8'b01100111: sig <= 8'b11001000;
            8'b01101000: sig <= 8'b11000101;
            8'b01101001: sig <= 8'b11000010;
            8'b01101010: sig <= 8'b11000000;
            8'b01101011: sig <= 8'b10111101;
            8'b01101100: sig <= 8'b10111010;
            8'b01101101: sig <= 8'b10111000;
            8'b01101110: sig <= 8'b10110101;
            8'b01101111: sig <= 8'b10110010;
            8'b01110000: sig <= 8'b10101111;
            8'b01110001: sig <= 8'b10101100;
            8'b01110010: sig <= 8'b10101001;
            8'b01110011: sig <= 8'b10100110;
            8'b01110100: sig <= 8'b10100011;
            8'b01110101: sig <= 8'b10100000;
            8'b01110110: sig <= 8'b10011101;
            8'b01110111: sig <= 8'b10011010;
            8'b01111000: sig <= 8'b10010111;
            8'b01111001: sig <= 8'b10010100;
            8'b01111010: sig <= 8'b10010001;
            8'b01111011: sig <= 8'b10001110;
            8'b01111100: sig <= 8'b10001011;
            8'b01111101: sig <= 8'b10001000;
            8'b01111110: sig <= 8'b10000101;
            8'b01111111: sig <= 8'b10000010;
            8'b10000000: sig <= 8'b01111111;
            8'b10000001: sig <= 8'b01111011;
            8'b10000010: sig <= 8'b01111000;
            8'b10000011: sig <= 8'b01110101;
            8'b10000100: sig <= 8'b01110010;
            8'b10000101: sig <= 8'b01101111;
            8'b10000110: sig <= 8'b01101100;
            8'b10000111: sig <= 8'b01101001;
            8'b10001000: sig <= 8'b01100110;
            8'b10001001: sig <= 8'b01100011;
            8'b10001010: sig <= 8'b01100000;
            8'b10001011: sig <= 8'b01011101;
            8'b10001100: sig <= 8'b01011010;
            8'b10001101: sig <= 8'b01010111;
            8'b10001110: sig <= 8'b01010100;
            8'b10001111: sig <= 8'b01010001;
            8'b10010000: sig <= 8'b01001110;
            8'b10010001: sig <= 8'b01001011;
            8'b10010010: sig <= 8'b01001000;
            8'b10010011: sig <= 8'b01000101;
            8'b10010100: sig <= 8'b01000011;
            8'b10010101: sig <= 8'b01000000;
            8'b10010110: sig <= 8'b00111101;
            8'b10010111: sig <= 8'b00111011;
            8'b10011000: sig <= 8'b00111000;
            8'b10011001: sig <= 8'b00110101;
            8'b10011010: sig <= 8'b00110011;
            8'b10011011: sig <= 8'b00110000;
            8'b10011100: sig <= 8'b00101110;
            8'b10011101: sig <= 8'b00101100;
            8'b10011110: sig <= 8'b00101001;
            8'b10011111: sig <= 8'b00100111;
            8'b10100000: sig <= 8'b00100101;
            8'b10100001: sig <= 8'b00100011;
            8'b10100010: sig <= 8'b00100000;
            8'b10100011: sig <= 8'b00011110;
            8'b10100100: sig <= 8'b00011100;
            8'b10100101: sig <= 8'b00011010;
            8'b10100110: sig <= 8'b00011000;
            8'b10100111: sig <= 8'b00010111;
            8'b10101000: sig <= 8'b00010101;
            8'b10101001: sig <= 8'b00010011;
            8'b10101010: sig <= 8'b00010010;
            8'b10101011: sig <= 8'b00010000;
            8'b10101100: sig <= 8'b00001110;
            8'b10101101: sig <= 8'b00001101;
            8'b10101110: sig <= 8'b00001100;
            8'b10101111: sig <= 8'b00001010;
            8'b10110000: sig <= 8'b00001001;
            8'b10110001: sig <= 8'b00001000;
            8'b10110010: sig <= 8'b00000111;
            8'b10110011: sig <= 8'b00000110;
            8'b10110100: sig <= 8'b00000101;
            8'b10110101: sig <= 8'b00000100;
            8'b10110110: sig <= 8'b00000011;
            8'b10110111: sig <= 8'b00000011;
            8'b10111000: sig <= 8'b00000010;
            8'b10111001: sig <= 8'b00000001;
            8'b10111010: sig <= 8'b00000001;
            8'b10111011: sig <= 8'b00000000;
            8'b10111100: sig <= 8'b00000000;
            8'b10111101: sig <= 8'b00000000;
            8'b10111110: sig <= 8'b00000000;
            8'b10111111: sig <= 8'b00000000;
            8'b11000000: sig <= 8'b00000000;
            8'b11000001: sig <= 8'b00000000;
            8'b11000010: sig <= 8'b00000000;
            8'b11000011: sig <= 8'b00000000;
            8'b11000100: sig <= 8'b00000000;
            8'b11000101: sig <= 8'b00000000;
            8'b11000110: sig <= 8'b00000001;
            8'b11000111: sig <= 8'b00000001;
            8'b11001000: sig <= 8'b00000010;
            8'b11001001: sig <= 8'b00000011;
            8'b11001010: sig <= 8'b00000011;
            8'b11001011: sig <= 8'b00000100;
            8'b11001100: sig <= 8'b00000101;
            8'b11001101: sig <= 8'b00000110;
            8'b11001110: sig <= 8'b00000111;
            8'b11001111: sig <= 8'b00001000;
            8'b11010000: sig <= 8'b00001001;
            8'b11010001: sig <= 8'b00001010;
            8'b11010010: sig <= 8'b00001100;
            8'b11010011: sig <= 8'b00001101;
            8'b11010100: sig <= 8'b00001110;
            8'b11010101: sig <= 8'b00010000;
            8'b11010110: sig <= 8'b00010010;
            8'b11010111: sig <= 8'b00010011;
            8'b11011000: sig <= 8'b00010101;
            8'b11011001: sig <= 8'b00010111;
            8'b11011010: sig <= 8'b00011000;
            8'b11011011: sig <= 8'b00011010;
            8'b11011100: sig <= 8'b00011100;
            8'b11011101: sig <= 8'b00011110;
            8'b11011110: sig <= 8'b00100000;
            8'b11011111: sig <= 8'b00100011;
            8'b11100000: sig <= 8'b00100101;
            8'b11100001: sig <= 8'b00100111;
            8'b11100010: sig <= 8'b00101001;
            8'b11100011: sig <= 8'b00101100;
            8'b11100100: sig <= 8'b00101110;
            8'b11100101: sig <= 8'b00110000;
            8'b11100110: sig <= 8'b00110011;
            8'b11100111: sig <= 8'b00110101;
            8'b11101000: sig <= 8'b00111000;
            8'b11101001: sig <= 8'b00111011;
            8'b11101010: sig <= 8'b00111101;
            8'b11101011: sig <= 8'b01000000;
            8'b11101100: sig <= 8'b01000011;
            8'b11101101: sig <= 8'b01000101;
            8'b11101110: sig <= 8'b01001000;
            8'b11101111: sig <= 8'b01001011;
            8'b11110000: sig <= 8'b01001110;
            8'b11110001: sig <= 8'b01010001;
            8'b11110010: sig <= 8'b01010100;
            8'b11110011: sig <= 8'b01010111;
            8'b11110100: sig <= 8'b01011010;
            8'b11110101: sig <= 8'b01011101;
            8'b11110110: sig <= 8'b01100000;
            8'b11110111: sig <= 8'b01100011;
            8'b11111000: sig <= 8'b01100110;
            8'b11111001: sig <= 8'b01101001;
            8'b11111010: sig <= 8'b01101100;
            8'b11111011: sig <= 8'b01101111;
            8'b11111100: sig <= 8'b01110010;
            8'b11111101: sig <= 8'b01110101;
            8'b11111110: sig <= 8'b01111000;
            8'b11111111: sig <= 8'b01111011;
            default: sig <= 8'b00000000; // should never happen
        endcase
    end
endmodule

